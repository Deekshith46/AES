module liner_tb;

reg
